--Library Declaration
library IEEE;
use IEEE.std_logic_1164.all;

package common is
   type matrix_type is array (natural range <>) of std_logic_vector (natural range <>);
end common;

package body common is
end common;
