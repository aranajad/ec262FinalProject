--Library Declaration
library IEEE;
use IEEE.std_logic_1164.all

--Entity Declaration
entity Register_64 is
    port (
        clk : in std_logic;
        rst : in std_logic;
        sig
    );
end Register_64;

architecture rtl of Register_64 is



begin



end architecture;